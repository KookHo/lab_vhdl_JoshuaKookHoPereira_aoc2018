library ieee;
use ieee.std_logic_1164.all;

entity portaAND is port(
	A: in STD_LOGIC;
	B: in STD_LOGIC;
	SA: out STD_LOGIC

);

end portaAND;

ARCHITECTURE behavior of portaAND is
BEGIN
	SA <= A and B;
END behavior;